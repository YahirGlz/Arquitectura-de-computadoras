module Jericalla(input [16:0], output reg [31:0]dataOut);

endmodule 